
`define	GPIO_CONFIG_ADDR        'd0
`define	GPIO_DOUT_ADDR          'd4
`define	GPIO_DIN_ADDR           'd8
`define	GPIO_DOUT_SET_ADDR      'd12
`define	GPIO_DOUT_CLR_ADDR      'd16

